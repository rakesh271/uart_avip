`ifndef UART_GLOBALS_PKG_INCLUDED_
`define UART_GLOBALS_PKG_INCLUDED_

//--------------------------------------------------------------------------------------------
// Package: uart_globals_pkg
// Used for storing enums, parameters and defines
//--------------------------------------------------------------------------------------------
package uart_globals_pkg;



endpackage: uart_globals_pkg

`endif
