//-------------------------------------------------------
//master monitor
//-------------------------------------------------------
module master_mon(uart_intf);

  initial
  begin
    $display("Master Monitor BFM");
  end

endmodule
