//-------------------------------------------------------
//master monitor bfm
//-------------------------------------------------------
module master_monitor_bfm(uart_if intf);

  initial
  begin
    $display("Master Monitor BFM");
  end

endmodule
